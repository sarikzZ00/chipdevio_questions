module multi_bit_fifo_tb;




initial begin
    $dumpfile("multi_bit_fifo.dump");
    $dumpvars( 0, multi_bit_fifo_tb_tb);
end

endmodule